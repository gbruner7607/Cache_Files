module way_arbiter #(
	parameter N_WAYS = 2,
	parameter AGE_WIDTH = 32
	)(

	);

endmodule : way_arbiter